module top_module (
    input clk,
    input slowena,
    input reset,
    output [3:0] q);
    
    always @(posedge clk) begin
        if (reset)
            q <= 4'h0;
        else if ((q == 4'h9) & slowena)
            q <= 4'h0;
        else if (slowena)
            q <= q + 1'b1;
    end

endmodule
